module pyramid_tb;

pyramid uut();
initial begin
        $display("start");
        $display("finish");

        $finish;

end
endmodule
