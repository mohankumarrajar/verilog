module reverse_pyramid_tb;
reverse_pyramid uut();

initial begin

        $display("start");
        $display("finish");

        $finish;
end
        endmodule
